
module Hazard_Unit(input  [4:0] Rs1D, Rs2D, Rs1E, Rs2E,
                input  [4:0] RdE, RdM, RdW,
                input  RegWriteM, RegWriteW,
					 input  ResultSrcE0, PCSrcE, rst,
                input  [31:0] InstrD,                      // Instruccion por ejecutar para saber cual pipeline
                output reg [1:0] ForwardAE, ForwardBE,      // Forward Pipeline Escalar
                output reg [1:0] VForwardAE, VForwardBE,    // Forward Pipeline Vectorial
                output StallD, StallF, FlushD, FlushE,      // Stalls y Flushes Escalares
                output VStallD, VStallF, VFlushD, VFlushE   // Stalls y Flushes Vectoriales
            );
					 


    wire lwStall;
    wire vLwStall;

    wire [6:0] funct7;
    wire [2:0] funct3;

    assign funct7 = InstrD[31:25];
    assign funct3 = InstrD[14:12];

    always @(*) begin
        ForwardAE = 2'b00;
        ForwardBE = 2'b00;
        VForwardAE = 2'b00;
        VForwardBE = 2'b00;

        if (funct7 == 7'b1010101) begin 
            if ((Rs1E == RdM) & (RegWriteM) & (Rs1E != 0)) // higher priority - most recent
                ForwardAE = 2'b10; // for forwarding ALU Result in Memory Stage
            else if ((Rs1E == RdW) & (RegWriteW) & (Rs1E != 0))
                ForwardAE = 2'b01; // for forwarding WriteBack Stage Result
                        
            if ((Rs2E == RdM) & (RegWriteM) & (Rs2E != 0))
                ForwardBE = 2'b10; // for forwarding ALU Result in Memory Stage
            else if ((Rs2E == RdW) & (RegWriteW) & (Rs2E != 0))
                ForwardBE = 2'b01; // for forwarding WriteBack Stage Result
        end else begin
            if ((Rs1E == RdM) & (RegWriteM) & (Rs1E != 0)) // higher priority - most recent
                VForwardAE = 2'b10; // for forwarding ALU Result in Memory Stage
            else if ((Rs1E == RdW) & (RegWriteW) & (Rs1E != 0))
                VForwardAE = 2'b01; // for forwarding WriteBack Stage Result
                        
            if ((Rs2E == RdM) & (RegWriteM) & (Rs2E != 0))
                VForwardBE = 2'b10; // for forwarding ALU Result in Memory Stage
            else if ((Rs2E == RdW) & (RegWriteW) & (Rs2E != 0))
                VForwardBE = 2'b01; // for forwarding WriteBack Stage Result
        end
    end


    assign lwStall = (ResultSrcE0 == 1) & ((RdE == Rs1D) | (RdE == Rs2D));
    assign vLwStall = (ResultSrcE0 == 1) & ((RdE == Rs1D) | (RdE == Rs2D));

    assign StallF = lwStall & (rst);
    assign StallD = lwStall & rst;
    assign FlushE = (lwStall | PCSrcE) & rst;
    assign FlushD = PCSrcE & rst;

    assign VStallF = vLwStall & (rst);
    assign VStallD = vLwStall & rst;
    assign VFlushE = (vLwStall | PCSrcE) & rst;
    assign VFlushD = PCSrcE & rst;


endmodule